`timescale 1ns/1ps

module ROM (addr,data);
input [31:0] addr;
output [31:0] data;

reg [31:0] data;
localparam ROM_size = 32;
reg [31:0] ROM_data[ROM_size-1:0];

always@(*)
	case(addr[8:2])	//addr : byte address -> addr[:2] word beginning address
		0: data <= 32'b00100100000000010000000000001000;
		1: data <= 32'b00110100000000100000000000000010;
		2: data <= 32'b00000000010000010001100000100000;
		3: data <= 32'b00000000011000100010100000100010;
		4: data <= 32'b00000000101000100010000000100100;
		5: data <= 32'b00000000100000100100000000100101;
		6: data <= 32'b00000000000010000100000001000000;
		7: data <= 32'b00010101000000011111111111111110;
		8: data <= 32'b00101000010001100000000000000100;
		9: data <= 32'b00101100110001110000000000000000;
		10: data <= 32'b00100100111001110000000000001000;
		11: data <= 32'b00010000111000011111111111111110;
		12: data <= 32'b10101100001000100000000000000100;
		13: data <= 32'b10001100001010010000000000000100;
		14: data <= 32'b00100101001010010000000000000000;
		15: data <= 32'b00100100000010101111111111111110;
		16: data <= 32'b00100101010010100000000000000001;
		17: data <= 32'b00110000010010110000000000000010;
		18: data <= 32'b00000000000000100101000000100001;
		19: data <= 32'b00000001010000100101000000100011;
		20: data <= 32'b00000001000000100101000000100110;
		21: data <= 32'b00000001000000100101000000100111;
		22: data <= 32'b00000001000000100101000000101011;
		23: data <= 32'b00000000000010000101000001000010;
		24: data <= 32'b00100000000010101111111111111111;
		25: data <= 32'b00000000000010100101100001000011;
		26: data <= 32'b11111100000000000000000000000000;
	   default:	data <= 32'h0000_0000;
	endcase
endmodule
